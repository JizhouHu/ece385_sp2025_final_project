module font_rom (
    input  logic [4:0] char_index,   // 0-23 
    input  logic [3:0] row,          // 0–15 for 8x16 font
    output logic [7:0] pixels        // 8 bits (left-to-right)
);

    logic [7:0] font [0:25][0:15];

    initial begin
        // --- T ---
        font[0][ 0] = 8'b00000000;
        font[0][ 1] = 8'b00000000;
        font[0][ 2] = 8'b11111111;
        font[0][ 3] = 8'b11011011;
        font[0][ 4] = 8'b10011001;
        font[0][ 5] = 8'b00011000;
        font[0][ 6] = 8'b00011000;
        font[0][ 7] = 8'b00011000;
        font[0][ 8] = 8'b00011000;
        font[0][ 9] = 8'b00011000;
        font[0][10] = 8'b00011000;
        font[0][11] = 8'b00111100;
        font[0][12] = 8'b00000000;
        font[0][13] = 8'b00000000;
        font[0][14] = 8'b00000000;
        font[0][15] = 8'b00000000;

        // --- A ---
        font[1][ 0] = 8'b00000000;
        font[1][ 1] = 8'b00000000;
        font[1][ 2] = 8'b00010000;
        font[1][ 3] = 8'b00111000;
        font[1][ 4] = 8'b01101100;
        font[1][ 5] = 8'b11000110;
        font[1][ 6] = 8'b11000110;
        font[1][ 7] = 8'b11111110;
        font[1][ 8] = 8'b11000110;
        font[1][ 9] = 8'b11000110;
        font[1][10] = 8'b11000110;
        font[1][11] = 8'b11000110;
        font[1][12] = 8'b00000000;
        font[1][13] = 8'b00000000;
        font[1][14] = 8'b00000000;
        font[1][15] = 8'b00000000;

        // --- N ---
        font[2][ 0] = 8'b00000000;
        font[2][ 1] = 8'b00000000;
        font[2][ 2] = 8'b11000110;
        font[2][ 3] = 8'b11100110;
        font[2][ 4] = 8'b11110110;
        font[2][ 5] = 8'b11111110;
        font[2][ 6] = 8'b11011110;
        font[2][ 7] = 8'b11001110;
        font[2][ 8] = 8'b11000110;
        font[2][ 9] = 8'b11000110;
        font[2][10] = 8'b11000110;
        font[2][11] = 8'b11000110;
        font[2][12] = 8'b00000000;
        font[2][13] = 8'b00000000;
        font[2][14] = 8'b00000000;
        font[2][15] = 8'b00000000;

        // --- K ---
        font[3][ 0] = 8'b00000000;
        font[3][ 1] = 8'b00000000;
        font[3][ 2] = 8'b11100110;
        font[3][ 3] = 8'b01100110;
        font[3][ 4] = 8'b01100110;
        font[3][ 5] = 8'b01101100;
        font[3][ 6] = 8'b01111000;
        font[3][ 7] = 8'b01111000;
        font[3][ 8] = 8'b01101100;
        font[3][ 9] = 8'b01100110;
        font[3][10] = 8'b01100110;
        font[3][11] = 8'b11100110;
        font[3][12] = 8'b00000000;
        font[3][13] = 8'b00000000;
        font[3][14] = 8'b00000000;
        font[3][15] = 8'b00000000;

        // --- 0 ---
        font[4][ 0] = 8'b00000000; // 0
        font[4][ 1] = 8'b00000000; // 1
        font[4][ 2] = 8'b01111100; // 2  *****
        font[4][ 3] = 8'b11000110; // 3 **   **
        font[4][ 4] = 8'b11000110; // 4 **   **
        font[4][ 5] = 8'b11001110; // 5 **  ***
        font[4][ 6] = 8'b11011110; // 6 ** ****
        font[4][ 7] = 8'b11110110; // 7 **** **
        font[4][ 8] = 8'b11100110; // 8 ***  **
        font[4][ 9] = 8'b11000110; // 9 **   **
        font[4][10] = 8'b11000110; // a **   **
        font[4][11] = 8'b01111100; // b  *****
        font[4][12] = 8'b00000000; // c
        font[4][13] = 8'b00000000; // d
        font[4][14] = 8'b00000000; // e
        font[4][15] = 8'b00000000; // f

        // --- W ---
        font[5][ 0] = 8'b00000000;
        font[5][ 1] = 8'b00000000;
        font[5][ 2] = 8'b11000011;
        font[5][ 3] = 8'b11000011;
        font[5][ 4] = 8'b11000011;
        font[5][ 5] = 8'b11000011;
        font[5][ 6] = 8'b11000011;
        font[5][ 7] = 8'b11011011;
        font[5][ 8] = 8'b11011011;
        font[5][ 9] = 8'b11111111;
        font[5][10] = 8'b01100110;
        font[5][11] = 8'b01100110;
        font[5][12] = 8'b00000000;
        font[5][13] = 8'b00000000;
        font[5][14] = 8'b00000000;
        font[5][15] = 8'b00000000;

        // --- R ---
        font[6][ 0] = 8'b00000000;
        font[6][ 1] = 8'b00000000;
        font[6][ 2] = 8'b11111100;
        font[6][ 3] = 8'b01100110;
        font[6][ 4] = 8'b01100110;
        font[6][ 5] = 8'b01100110;
        font[6][ 6] = 8'b01111100;
        font[6][ 7] = 8'b01101100;
        font[6][ 8] = 8'b01100110;
        font[6][ 9] = 8'b01100110;
        font[6][10] = 8'b01100110;
        font[6][11] = 8'b11100110;
        font[6][12] = 8'b00000000;
        font[6][13] = 8'b00000000;
        font[6][14] = 8'b00000000;
        font[6][15] = 8'b00000000;

        // --- B ---
        font[7][ 0] = 8'b00000000; //                    
        font[7][ 1] = 8'b00000000; //                    
        font[7][ 2] = 8'b11111100; // ******            
        font[7][ 3] = 8'b01100110; //  **  **           
        font[7][ 4] = 8'b01100110; //  **  **           
        font[7][ 5] = 8'b01100110; //  **  **           
        font[7][ 6] = 8'b01111100; //  *****            
        font[7][ 7] = 8'b01100110; //  **  **           
        font[7][ 8] = 8'b01100110; //  **  **           
        font[7][ 9] = 8'b01100110; //  **  **           
        font[7][10] = 8'b01100110; //  **  **           
        font[7][11] = 8'b11111100; // ******            
        font[7][12] = 8'b00000000; //                    
        font[7][13] = 8'b00000000; //                    
        font[7][14] = 8'b00000000; //                    
        font[7][15] = 8'b00000000; //    

        // --- P ---
        font[8][ 0] = 8'b00000000; // 0
        font[8][ 1] = 8'b00000000; // 1
        font[8][ 2] = 8'b11111100; // 2 ******
        font[8][ 3] = 8'b01100110; // 3  **  **
        font[8][ 4] = 8'b01100110; // 4  **  **
        font[8][ 5] = 8'b01100110; // 5  **  **
        font[8][ 6] = 8'b01111100; // 6  *****
        font[8][ 7] = 8'b01100000; // 7  **
        font[8][ 8] = 8'b01100000; // 8  **
        font[8][ 9] = 8'b01100000; // 9  **
        font[8][10] = 8'b01100000; // a  **
        font[8][11] = 8'b11110000; // b ****
        font[8][12] = 8'b00000000; // c
        font[8][13] = 8'b00000000; // d
        font[8][14] = 8'b00000000; // e
        font[8][15] = 8'b00000000; // f

        // --- E ---
        font[9][ 0] = 8'b00000000; // 0
        font[9][ 1] = 8'b00000000; // 1
        font[9][ 2] = 8'b11111110; // 2 *******
        font[9][ 3] = 8'b01100110; // 3  **  **
        font[9][ 4] = 8'b01100010; // 4  **   *
        font[9][ 5] = 8'b01101000; // 5  ** *
        font[9][ 6] = 8'b01111000; // 6  ****
        font[9][ 7] = 8'b01101000; // 7  ** *
        font[9][ 8] = 8'b01100000; // 8  **
        font[9][ 9] = 8'b01100010; // 9  **   *
        font[9][10] = 8'b01100110; // a  **  **
        font[9][11] = 8'b11111110; // b *******
        font[9][12] = 8'b00000000; // c
        font[9][13] = 8'b00000000; // d
        font[9][14] = 8'b00000000; // e
        font[9][15] = 8'b00000000; // f

        // --- F ---
        font[10][ 0] = 8'b00000000; // 0
        font[10][ 1] = 8'b00000000; // 1
        font[10][ 2] = 8'b11111110; // 2 *******
        font[10][ 3] = 8'b01100110; // 3  **  **
        font[10][ 4] = 8'b01100010; // 4  **   *
        font[10][ 5] = 8'b01101000; // 5  ** *
        font[10][ 6] = 8'b01111000; // 6  ****
        font[10][ 7] = 8'b01101000; // 7  ** *
        font[10][ 8] = 8'b01100000; // 8  **
        font[10][ 9] = 8'b01100000; // 9  **
        font[10][10] = 8'b01100000; // a  **
        font[10][11] = 8'b11110000; // b ****
        font[10][12] = 8'b00000000; // c
        font[10][13] = 8'b00000000; // d
        font[10][14] = 8'b00000000; // e
        font[10][15] = 8'b00000000; // f

        // --- I ---
        font[11][ 0] = 8'b00000000; // 0
        font[11][ 1] = 8'b00000000; // 1
        font[11][ 2] = 8'b00111100; // 2   ****
        font[11][ 3] = 8'b00011000; // 3    **
        font[11][ 4] = 8'b00011000; // 4    **
        font[11][ 5] = 8'b00011000; // 5    **
        font[11][ 6] = 8'b00011000; // 6    **
        font[11][ 7] = 8'b00011000; // 7    **
        font[11][ 8] = 8'b00011000; // 8    **
        font[11][ 9] = 8'b00011000; // 9    **
        font[11][10] = 8'b00011000; // a    **
        font[11][11] = 8'b00111100; // b   ****
        font[11][12] = 8'b00000000; // c
        font[11][13] = 8'b00000000; // d
        font[11][14] = 8'b00000000; // e
        font[11][15] = 8'b00000000; // f

        // --- L ---
        font[12][ 0] = 8'b00000000; // 0
        font[12][ 1] = 8'b00000000; // 1
        font[12][ 2] = 8'b11110000; // 2 ****
        font[12][ 3] = 8'b01100000; // 3  **
        font[12][ 4] = 8'b01100000; // 4  **
        font[12][ 5] = 8'b01100000; // 5  **
        font[12][ 6] = 8'b01100000; // 6  **
        font[12][ 7] = 8'b01100000; // 7  **
        font[12][ 8] = 8'b01100000; // 8  **
        font[12][ 9] = 8'b01100010; // 9  **   *
        font[12][10] = 8'b01100110; // a  **  **
        font[12][11] = 8'b11111110; // b *******
        font[12][12] = 8'b00000000; // c
        font[12][13] = 8'b00000000; // d
        font[12][14] = 8'b00000000; // e
        font[12][15] = 8'b00000000; // f

        // error position (originally store M) M: 24
        // might read wrong pixels from error position
        font[13][ 0] = 8'b00000000; // 0
        font[13][ 1] = 8'b00000000; // 1
        font[13][ 2] = 8'b11000011; // 2 **    **
        font[13][ 3] = 8'b11100111; // 3 ***  ***
        font[13][ 4] = 8'b11111111; // 4 ********
        font[13][ 5] = 8'b11111111; // 5 ********
        font[13][ 6] = 8'b11011011; // 6 ** ** **
        font[13][ 7] = 8'b11000011; // 7 **    **
        font[13][ 8] = 8'b11000011; // 8 **    **
        font[13][ 9] = 8'b11000011; // 9 **    **
        font[13][10] = 8'b11000011; // a **    **
        font[13][11] = 8'b11000011; // b **    **
        font[13][12] = 8'b00000000; // c
        font[13][13] = 8'b00000000; // d
        font[13][14] = 8'b00000000; // e
        font[13][15] = 8'b00000000; // f

        // error position (originally store 0) 0: 4
        font[14][ 0] = 8'b00000000; // 0
        font[14][ 1] = 8'b00000000; // 1
        font[14][ 2] = 8'b01111100; // 2  *****
        font[14][ 3] = 8'b11000110; // 3 **   **
        font[14][ 4] = 8'b11000110; // 4 **   **
        font[13][ 5] = 8'b11001110; // 5 **  ***
        font[14][ 6] = 8'b11011110; // 6 ** ****
        font[14][ 7] = 8'b11110110; // 7 **** **
        font[14][ 8] = 8'b11100110; // 8 ***  **
        font[14][ 9] = 8'b11000110; // 9 **   **
        font[14][10] = 8'b11000110; // a **   **
        font[14][11] = 8'b01111100; // b  *****
        font[14][12] = 8'b00000000; // c
        font[14][13] = 8'b00000000; // d
        font[14][14] = 8'b00000000; // e
        font[14][15] = 8'b00000000; // f
        
        // --- 1 ---
        font[15][ 0] = 8'b00000000; // 0
        font[15][ 1] = 8'b00000000; // 1
        font[15][ 2] = 8'b00011000; // 2
        font[15][ 3] = 8'b00111000; // 3
        font[15][ 4] = 8'b01111000; // 4    **
        font[15][ 5] = 8'b00011000; // 5   ***
        font[15][ 6] = 8'b00011000; // 6  ****
        font[15][ 7] = 8'b00011000; // 7    **
        font[15][ 8] = 8'b00011000; // 8    **
        font[15][ 9] = 8'b00011000; // 9    **
        font[15][10] = 8'b00011000; // a    **
        font[15][11] = 8'b01111110; // b    **
        font[15][12] = 8'b00000000; // c    **
        font[15][13] = 8'b00000000; // d  ******
        font[15][14] = 8'b00000000; // e
        font[15][15] = 8'b00000000; // f

         // --- 2 ---
        font[16][ 0] = 8'b00000000;
        font[16][ 1] = 8'b00000000;
        font[16][ 2] = 8'b01111100; //  *****
        font[16][ 3] = 8'b11000110; // **   **
        font[16][ 4] = 8'b00000110; //      **
        font[16][ 5] = 8'b00001100; //     **
        font[16][ 6] = 8'b00011000; //    **
        font[16][ 7] = 8'b00110000; //   **
        font[16][ 8] = 8'b01100000; //  **
        font[16][ 9] = 8'b11000000; // **
        font[16][10] = 8'b11000110; // **   **
        font[16][11] = 8'b11111110; // *******
        font[16][12] = 8'b00000000;
        font[16][13] = 8'b00000000;
        font[16][14] = 8'b00000000;
        font[16][15] = 8'b00000000;
        
        // --- 3 ---
        font[17][ 0] = 8'b00000000;
        font[17][ 1] = 8'b00000000;
        font[17][ 2] = 8'b01111100; //  *****
        font[17][ 3] = 8'b11000110; // **   **
        font[17][ 4] = 8'b00000110; //      **
        font[17][ 5] = 8'b00000110; //      **
        font[17][ 6] = 8'b00111100; //   ****
        font[17][ 7] = 8'b00000110; //      **
        font[17][ 8] = 8'b00000110; //      **
        font[17][ 9] = 8'b00000110; //      **
        font[17][10] = 8'b11000110; // **   **
        font[17][11] = 8'b01111100; //  *****
        font[17][12] = 8'b00000000;
        font[17][13] = 8'b00000000;
        font[17][14] = 8'b00000000;
        font[17][15] = 8'b00000000;
         
        // --- 4 ---
        font[18][ 0] = 8'b00000000;
        font[18][ 1] = 8'b00000000;
        font[18][ 2] = 8'b00001100; //     **
        font[18][ 3] = 8'b00011100; //    ***
        font[18][ 4] = 8'b00111100; //   ****
        font[18][ 5] = 8'b01101100; //  ** **
        font[18][ 6] = 8'b11001100; // **  **
        font[18][ 7] = 8'b11111110; // *******
        font[18][ 8] = 8'b00001100; //     **
        font[18][ 9] = 8'b00001100; //     **
        font[18][10] = 8'b00001100; //     **
        font[18][11] = 8'b00011110; //    ****
        font[18][12] = 8'b00000000;
        font[18][13] = 8'b00000000;
        font[18][14] = 8'b00000000;
        font[18][15] = 8'b00000000;

        // --- 5 ---
        font[19][ 0] = 8'b00000000;
        font[19][ 1] = 8'b00000000;
        font[19][ 2] = 8'b11111110; // *******
        font[19][ 3] = 8'b11000000; // **
        font[19][ 4] = 8'b11000000; // **
        font[19][ 5] = 8'b11000000; // **
        font[19][ 6] = 8'b11111100; // ******
        font[19][ 7] = 8'b00000110; //      **
        font[19][ 8] = 8'b00000110; //      **
        font[19][ 9] = 8'b00000110; //      **
        font[19][10] = 8'b11000110; // **   **
        font[19][11] = 8'b01111100; //  *****
        font[19][12] = 8'b00000000;
        font[19][13] = 8'b00000000;
        font[19][14] = 8'b00000000;
        font[19][15] = 8'b00000000;

        // --- 6 ---
        font[20][ 0] = 8'b00000000;
        font[20][ 1] = 8'b00000000;
        font[20][ 2] = 8'b00111000; //   ***
        font[20][ 3] = 8'b01100000; //  **
        font[20][ 4] = 8'b11000000; // **
        font[20][ 5] = 8'b11000000; // **
        font[20][ 6] = 8'b11111100; // ******
        font[20][ 7] = 8'b11000110; // **   **
        font[20][ 8] = 8'b11000110; // **   **
        font[20][ 9] = 8'b11000110; // **   **
        font[20][10] = 8'b11000110; // **   **
        font[20][11] = 8'b01111100; //  *****
        font[20][12] = 8'b00000000;
        font[20][13] = 8'b00000000;
        font[20][14] = 8'b00000000;
        font[20][15] = 8'b00000000;

        // --- 7 ---
        font[21][ 0] = 8'b00000000;
        font[21][ 1] = 8'b00000000;
        font[21][ 2] = 8'b11111110; // *******
        font[21][ 3] = 8'b11000110; // **   **
        font[21][ 4] = 8'b00000110; //      **
        font[21][ 5] = 8'b00000110; //      **
        font[21][ 6] = 8'b00001100; //     **
        font[21][ 7] = 8'b00011000; //    **
        font[21][ 8] = 8'b00110000; //   **
        font[21][ 9] = 8'b00110000; //   **
        font[21][10] = 8'b00110000; //   **
        font[21][11] = 8'b00110000; //   **
        font[21][12] = 8'b00000000;
        font[21][13] = 8'b00000000;
        font[21][14] = 8'b00000000;
        font[21][15] = 8'b00000000;
        
        // --- 8 ---
        font[22][ 0] = 8'b00000000;
        font[22][ 1] = 8'b00000000;
        font[22][ 2] = 8'b01111100; //  *****
        font[22][ 3] = 8'b11000110; // **   **
        font[22][ 4] = 8'b11000110; // **   **
        font[22][ 5] = 8'b11000110; // **   **
        font[22][ 6] = 8'b01111100; //  *****
        font[22][ 7] = 8'b11000110; // **   **
        font[22][ 8] = 8'b11000110; // **   **
        font[22][ 9] = 8'b11000110; // **   **
        font[22][10] = 8'b11000110; // **   **
        font[22][11] = 8'b01111100; //  *****
        font[22][12] = 8'b00000000;
        font[22][13] = 8'b00000000;
        font[22][14] = 8'b00000000;
        font[22][15] = 8'b00000000;
    
        // --- 9 ---
        font[23][ 0] = 8'b00000000;
        font[23][ 1] = 8'b00000000;
        font[23][ 2] = 8'b01111100; //  *****
        font[23][ 3] = 8'b11000110; // **   **
        font[23][ 4] = 8'b11000110; // **   **
        font[23][ 5] = 8'b11000110; // **   **
        font[23][ 6] = 8'b01111110; //  ******
        font[23][ 7] = 8'b00000110; //      **
        font[23][ 8] = 8'b00000110; //      **
        font[23][ 9] = 8'b00000110; //      **
        font[23][10] = 8'b00001100; //     **
        font[23][11] = 8'b01111000; //  ****
        font[23][12] = 8'b00000000;
        font[23][13] = 8'b00000000;
        font[23][14] = 8'b00000000;
        font[23][15] = 8'b00000000;

        // --- M ---
        font[24][ 0] = 8'b00000000; // 0
        font[24][ 1] = 8'b00000000; // 1
        font[24][ 2] = 8'b11000011; // 2 **    **
        font[24][ 3] = 8'b11100111; // 3 ***  ***
        font[24][ 4] = 8'b11111111; // 4 ********
        font[24][ 5] = 8'b11111111; // 5 ********
        font[24][ 6] = 8'b11011011; // 6 ** ** **
        font[24][ 7] = 8'b11000011; // 7 **    **
        font[24][ 8] = 8'b11000011; // 8 **    **
        font[24][ 9] = 8'b11000011; // 9 **    **
        font[24][10] = 8'b11000011; // a **    **
        font[24][11] = 8'b11000011; // b **    **
        font[24][12] = 8'b00000000; // c
        font[24][13] = 8'b00000000; // d
        font[24][14] = 8'b00000000; // e
        font[24][15] = 8'b00000000; // f

        // --- Space --- (space can be store in "error" position)
        font[25][ 0] = 8'b00000000;
        font[25][ 1] = 8'b00000000;
        font[25][ 2] = 8'b00000000;
        font[25][ 3] = 8'b00000000;
        font[25][ 4] = 8'b00000000;
        font[25][ 5] = 8'b00000000;
        font[25][ 6] = 8'b00000000;
        font[25][ 7] = 8'b00000000;
        font[25][ 8] = 8'b00000000;
        font[25][ 9] = 8'b00000000;
        font[25][10] = 8'b00000000;
        font[25][11] = 8'b00000000;
        font[25][12] = 8'b00000000;
        font[25][13] = 8'b00000000;
        font[25][14] = 8'b00000000;
        font[25][15] = 8'b00000000;
    end

    // Output the row
    assign pixels = font[char_index][row];

endmodule
         